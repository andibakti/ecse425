library ieee;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity id_reg is 
	port(
		cl
		);

end id_reg;
